// olive_std_core.v

// Generated using ACDS version 17.0 602

`timescale 1 ps / 1 ps
module olive_std_core (
		input  wire        clk_100m_clk,           // clk_100m.clk
		input  wire        clk_25m_clk,            //  clk_25m.clk
		output wire        epcs_ss_n,              //     epcs.ss_n
		output wire        epcs_sclk,              //         .sclk
		output wire        epcs_mosi,              //         .mosi
		input  wire        epcs_miso,              //         .miso
		input  wire        hostuart_rxd,           // hostuart.rxd
		output wire        hostuart_txd,           //         .txd
		input  wire        i2c_scl,                //      i2c.scl
		output wire        i2c_scl_oe,             //         .scl_oe
		input  wire        i2c_sda,                //         .sda
		output wire        i2c_sda_oe,             //         .sda_oe
		output wire        led_export,             //      led.export
		input  wire        nios2_cpu_resetrequest, //    nios2.cpu_resetrequest
		output wire        nios2_cpu_resettaken,   //         .cpu_resettaken
		output wire        pfcif_pfc_clk,          //    pfcif.pfc_clk
		output wire        pfcif_pfc_reset,        //         .pfc_reset
		output wire [36:0] pfcif_cmd,              //         .cmd
		input  wire [31:0] pfcif_resp,             //         .resp
		input  wire        reset_reset_n,          //    reset.reset_n
		output wire [11:0] sdr_addr,               //      sdr.addr
		output wire [1:0]  sdr_ba,                 //         .ba
		output wire        sdr_cas_n,              //         .cas_n
		output wire        sdr_cke,                //         .cke
		output wire        sdr_cs_n,               //         .cs_n
		inout  wire [15:0] sdr_dq,                 //         .dq
		output wire [1:0]  sdr_dqm,                //         .dqm
		output wire        sdr_ras_n,              //         .ras_n
		output wire        sdr_we_n,               //         .we_n
		output wire [7:0]  servo_pwm,              //    servo.pwm
		output wire [7:0]  servo_dsm,              //         .dsm
		output wire        spi_ss_n,               //      spi.ss_n
		output wire        spi_sclk,               //         .sclk
		output wire        spi_mosi,               //         .mosi
		input  wire        spi_miso,               //         .miso
		input  wire        uart0_rxd,              //    uart0.rxd
		output wire        uart0_txd,              //         .txd
		input  wire        uart0_cts_n,            //         .cts_n
		output wire        uart0_rts_n,            //         .rts_n
		input  wire        uart1_rxd,              //    uart1.rxd
		output wire        uart1_txd,              //         .txd
		input  wire        uart1_cts_n,            //         .cts_n
		output wire        uart1_rts_n             //         .rts_n
	);

	wire  [31:0] nios2_fast_data_master_readdata;                          // mm_interconnect_0:nios2_fast_data_master_readdata -> nios2_fast:d_readdata
	wire         nios2_fast_data_master_waitrequest;                       // mm_interconnect_0:nios2_fast_data_master_waitrequest -> nios2_fast:d_waitrequest
	wire         nios2_fast_data_master_debugaccess;                       // nios2_fast:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_fast_data_master_debugaccess
	wire  [28:0] nios2_fast_data_master_address;                           // nios2_fast:d_address -> mm_interconnect_0:nios2_fast_data_master_address
	wire   [3:0] nios2_fast_data_master_byteenable;                        // nios2_fast:d_byteenable -> mm_interconnect_0:nios2_fast_data_master_byteenable
	wire         nios2_fast_data_master_read;                              // nios2_fast:d_read -> mm_interconnect_0:nios2_fast_data_master_read
	wire         nios2_fast_data_master_readdatavalid;                     // mm_interconnect_0:nios2_fast_data_master_readdatavalid -> nios2_fast:d_readdatavalid
	wire         nios2_fast_data_master_write;                             // nios2_fast:d_write -> mm_interconnect_0:nios2_fast_data_master_write
	wire  [31:0] nios2_fast_data_master_writedata;                         // nios2_fast:d_writedata -> mm_interconnect_0:nios2_fast_data_master_writedata
	wire  [31:0] nios2_fast_instruction_master_readdata;                   // mm_interconnect_0:nios2_fast_instruction_master_readdata -> nios2_fast:i_readdata
	wire         nios2_fast_instruction_master_waitrequest;                // mm_interconnect_0:nios2_fast_instruction_master_waitrequest -> nios2_fast:i_waitrequest
	wire  [27:0] nios2_fast_instruction_master_address;                    // nios2_fast:i_address -> mm_interconnect_0:nios2_fast_instruction_master_address
	wire         nios2_fast_instruction_master_read;                       // nios2_fast:i_read -> mm_interconnect_0:nios2_fast_instruction_master_read
	wire         nios2_fast_instruction_master_readdatavalid;              // mm_interconnect_0:nios2_fast_instruction_master_readdatavalid -> nios2_fast:i_readdatavalid
	wire  [31:0] mm_interconnect_0_ufm_data_readdata;                      // ufm:avmm_data_readdata -> mm_interconnect_0:ufm_data_readdata
	wire         mm_interconnect_0_ufm_data_waitrequest;                   // ufm:avmm_data_waitrequest -> mm_interconnect_0:ufm_data_waitrequest
	wire  [12:0] mm_interconnect_0_ufm_data_address;                       // mm_interconnect_0:ufm_data_address -> ufm:avmm_data_addr
	wire         mm_interconnect_0_ufm_data_read;                          // mm_interconnect_0:ufm_data_read -> ufm:avmm_data_read
	wire         mm_interconnect_0_ufm_data_readdatavalid;                 // ufm:avmm_data_readdatavalid -> mm_interconnect_0:ufm_data_readdatavalid
	wire   [1:0] mm_interconnect_0_ufm_data_burstcount;                    // mm_interconnect_0:ufm_data_burstcount -> ufm:avmm_data_burstcount
	wire  [31:0] mm_interconnect_0_nios2_fast_debug_mem_slave_readdata;    // nios2_fast:debug_mem_slave_readdata -> mm_interconnect_0:nios2_fast_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_fast_debug_mem_slave_waitrequest; // nios2_fast:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_fast_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_fast_debug_mem_slave_debugaccess; // mm_interconnect_0:nios2_fast_debug_mem_slave_debugaccess -> nios2_fast:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_fast_debug_mem_slave_address;     // mm_interconnect_0:nios2_fast_debug_mem_slave_address -> nios2_fast:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_fast_debug_mem_slave_read;        // mm_interconnect_0:nios2_fast_debug_mem_slave_read -> nios2_fast:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_fast_debug_mem_slave_byteenable;  // mm_interconnect_0:nios2_fast_debug_mem_slave_byteenable -> nios2_fast:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_fast_debug_mem_slave_write;       // mm_interconnect_0:nios2_fast_debug_mem_slave_write -> nios2_fast:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_fast_debug_mem_slave_writedata;   // mm_interconnect_0:nios2_fast_debug_mem_slave_writedata -> nios2_fast:debug_mem_slave_writedata
	wire  [31:0] mm_interconnect_0_peripheral_bridge_s0_readdata;          // peripheral_bridge:s0_readdata -> mm_interconnect_0:peripheral_bridge_s0_readdata
	wire         mm_interconnect_0_peripheral_bridge_s0_waitrequest;       // peripheral_bridge:s0_waitrequest -> mm_interconnect_0:peripheral_bridge_s0_waitrequest
	wire         mm_interconnect_0_peripheral_bridge_s0_debugaccess;       // mm_interconnect_0:peripheral_bridge_s0_debugaccess -> peripheral_bridge:s0_debugaccess
	wire   [8:0] mm_interconnect_0_peripheral_bridge_s0_address;           // mm_interconnect_0:peripheral_bridge_s0_address -> peripheral_bridge:s0_address
	wire         mm_interconnect_0_peripheral_bridge_s0_read;              // mm_interconnect_0:peripheral_bridge_s0_read -> peripheral_bridge:s0_read
	wire   [3:0] mm_interconnect_0_peripheral_bridge_s0_byteenable;        // mm_interconnect_0:peripheral_bridge_s0_byteenable -> peripheral_bridge:s0_byteenable
	wire         mm_interconnect_0_peripheral_bridge_s0_readdatavalid;     // peripheral_bridge:s0_readdatavalid -> mm_interconnect_0:peripheral_bridge_s0_readdatavalid
	wire         mm_interconnect_0_peripheral_bridge_s0_write;             // mm_interconnect_0:peripheral_bridge_s0_write -> peripheral_bridge:s0_write
	wire  [31:0] mm_interconnect_0_peripheral_bridge_s0_writedata;         // mm_interconnect_0:peripheral_bridge_s0_writedata -> peripheral_bridge:s0_writedata
	wire   [0:0] mm_interconnect_0_peripheral_bridge_s0_burstcount;        // mm_interconnect_0:peripheral_bridge_s0_burstcount -> peripheral_bridge:s0_burstcount
	wire         mm_interconnect_0_sdram_s1_chipselect;                    // mm_interconnect_0:sdram_s1_chipselect -> sdram:az_cs
	wire  [15:0] mm_interconnect_0_sdram_s1_readdata;                      // sdram:za_data -> mm_interconnect_0:sdram_s1_readdata
	wire         mm_interconnect_0_sdram_s1_waitrequest;                   // sdram:za_waitrequest -> mm_interconnect_0:sdram_s1_waitrequest
	wire  [21:0] mm_interconnect_0_sdram_s1_address;                       // mm_interconnect_0:sdram_s1_address -> sdram:az_addr
	wire         mm_interconnect_0_sdram_s1_read;                          // mm_interconnect_0:sdram_s1_read -> sdram:az_rd_n
	wire   [1:0] mm_interconnect_0_sdram_s1_byteenable;                    // mm_interconnect_0:sdram_s1_byteenable -> sdram:az_be_n
	wire         mm_interconnect_0_sdram_s1_readdatavalid;                 // sdram:za_valid -> mm_interconnect_0:sdram_s1_readdatavalid
	wire         mm_interconnect_0_sdram_s1_write;                         // mm_interconnect_0:sdram_s1_write -> sdram:az_wr_n
	wire  [15:0] mm_interconnect_0_sdram_s1_writedata;                     // mm_interconnect_0:sdram_s1_writedata -> sdram:az_data
	wire  [31:0] mm_interconnect_0_epcs_s1_readdata;                       // epcs:avs_readdata -> mm_interconnect_0:epcs_s1_readdata
	wire   [0:0] mm_interconnect_0_epcs_s1_address;                        // mm_interconnect_0:epcs_s1_address -> epcs:avs_address
	wire         mm_interconnect_0_epcs_s1_read;                           // mm_interconnect_0:epcs_s1_read -> epcs:avs_read
	wire         mm_interconnect_0_epcs_s1_write;                          // mm_interconnect_0:epcs_s1_write -> epcs:avs_write
	wire  [31:0] mm_interconnect_0_epcs_s1_writedata;                      // mm_interconnect_0:epcs_s1_writedata -> epcs:avs_writedata
	wire         peripheral_bridge_m0_waitrequest;                         // mm_interconnect_1:peripheral_bridge_m0_waitrequest -> peripheral_bridge:m0_waitrequest
	wire  [31:0] peripheral_bridge_m0_readdata;                            // mm_interconnect_1:peripheral_bridge_m0_readdata -> peripheral_bridge:m0_readdata
	wire         peripheral_bridge_m0_debugaccess;                         // peripheral_bridge:m0_debugaccess -> mm_interconnect_1:peripheral_bridge_m0_debugaccess
	wire   [8:0] peripheral_bridge_m0_address;                             // peripheral_bridge:m0_address -> mm_interconnect_1:peripheral_bridge_m0_address
	wire         peripheral_bridge_m0_read;                                // peripheral_bridge:m0_read -> mm_interconnect_1:peripheral_bridge_m0_read
	wire   [3:0] peripheral_bridge_m0_byteenable;                          // peripheral_bridge:m0_byteenable -> mm_interconnect_1:peripheral_bridge_m0_byteenable
	wire         peripheral_bridge_m0_readdatavalid;                       // mm_interconnect_1:peripheral_bridge_m0_readdatavalid -> peripheral_bridge:m0_readdatavalid
	wire  [31:0] peripheral_bridge_m0_writedata;                           // peripheral_bridge:m0_writedata -> mm_interconnect_1:peripheral_bridge_m0_writedata
	wire         peripheral_bridge_m0_write;                               // peripheral_bridge:m0_write -> mm_interconnect_1:peripheral_bridge_m0_write
	wire   [0:0] peripheral_bridge_m0_burstcount;                          // peripheral_bridge:m0_burstcount -> mm_interconnect_1:peripheral_bridge_m0_burstcount
	wire  [31:0] mm_interconnect_1_dual_boot_0_avalon_readdata;            // dual_boot_0:avmm_rcv_readdata -> mm_interconnect_1:dual_boot_0_avalon_readdata
	wire   [2:0] mm_interconnect_1_dual_boot_0_avalon_address;             // mm_interconnect_1:dual_boot_0_avalon_address -> dual_boot_0:avmm_rcv_address
	wire         mm_interconnect_1_dual_boot_0_avalon_read;                // mm_interconnect_1:dual_boot_0_avalon_read -> dual_boot_0:avmm_rcv_read
	wire         mm_interconnect_1_dual_boot_0_avalon_write;               // mm_interconnect_1:dual_boot_0_avalon_write -> dual_boot_0:avmm_rcv_write
	wire  [31:0] mm_interconnect_1_dual_boot_0_avalon_writedata;           // mm_interconnect_1:dual_boot_0_avalon_writedata -> dual_boot_0:avmm_rcv_writedata
	wire  [31:0] mm_interconnect_1_pfc_avalon_slave_readdata;              // pfc:avs_readdata -> mm_interconnect_1:pfc_avalon_slave_readdata
	wire   [3:0] mm_interconnect_1_pfc_avalon_slave_address;               // mm_interconnect_1:pfc_avalon_slave_address -> pfc:avs_address
	wire         mm_interconnect_1_pfc_avalon_slave_read;                  // mm_interconnect_1:pfc_avalon_slave_read -> pfc:avs_read
	wire         mm_interconnect_1_pfc_avalon_slave_write;                 // mm_interconnect_1:pfc_avalon_slave_write -> pfc:avs_write
	wire  [31:0] mm_interconnect_1_pfc_avalon_slave_writedata;             // mm_interconnect_1:pfc_avalon_slave_writedata -> pfc:avs_writedata
	wire  [31:0] mm_interconnect_1_servo_avalon_slave_readdata;            // servo:avs_readdata -> mm_interconnect_1:servo_avalon_slave_readdata
	wire   [4:0] mm_interconnect_1_servo_avalon_slave_address;             // mm_interconnect_1:servo_avalon_slave_address -> servo:avs_address
	wire         mm_interconnect_1_servo_avalon_slave_read;                // mm_interconnect_1:servo_avalon_slave_read -> servo:avs_read
	wire         mm_interconnect_1_servo_avalon_slave_write;               // mm_interconnect_1:servo_avalon_slave_write -> servo:avs_write
	wire  [31:0] mm_interconnect_1_servo_avalon_slave_writedata;           // mm_interconnect_1:servo_avalon_slave_writedata -> servo:avs_writedata
	wire  [31:0] mm_interconnect_1_chipid_chipid_readdata;                 // chipid:chipid_readdata -> mm_interconnect_1:chipid_chipid_readdata
	wire         mm_interconnect_1_chipid_chipid_waitrequest;              // chipid:chipid_waitrequest -> mm_interconnect_1:chipid_chipid_waitrequest
	wire   [0:0] mm_interconnect_1_chipid_chipid_address;                  // mm_interconnect_1:chipid_chipid_address -> chipid:chipid_address
	wire         mm_interconnect_1_chipid_chipid_read;                     // mm_interconnect_1:chipid_chipid_read -> chipid:chipid_read
	wire  [31:0] mm_interconnect_1_sysid_control_slave_readdata;           // sysid:readdata -> mm_interconnect_1:sysid_control_slave_readdata
	wire   [0:0] mm_interconnect_1_sysid_control_slave_address;            // mm_interconnect_1:sysid_control_slave_address -> sysid:address
	wire         mm_interconnect_1_systimer_s1_chipselect;                 // mm_interconnect_1:systimer_s1_chipselect -> systimer:chipselect
	wire  [15:0] mm_interconnect_1_systimer_s1_readdata;                   // systimer:readdata -> mm_interconnect_1:systimer_s1_readdata
	wire   [2:0] mm_interconnect_1_systimer_s1_address;                    // mm_interconnect_1:systimer_s1_address -> systimer:address
	wire         mm_interconnect_1_systimer_s1_write;                      // mm_interconnect_1:systimer_s1_write -> systimer:write_n
	wire  [15:0] mm_interconnect_1_systimer_s1_writedata;                  // mm_interconnect_1:systimer_s1_writedata -> systimer:writedata
	wire         mm_interconnect_1_uart0_s1_chipselect;                    // mm_interconnect_1:uart0_s1_chipselect -> uart0:chipselect
	wire  [15:0] mm_interconnect_1_uart0_s1_readdata;                      // uart0:readdata -> mm_interconnect_1:uart0_s1_readdata
	wire   [2:0] mm_interconnect_1_uart0_s1_address;                       // mm_interconnect_1:uart0_s1_address -> uart0:address
	wire         mm_interconnect_1_uart0_s1_read;                          // mm_interconnect_1:uart0_s1_read -> uart0:read_n
	wire         mm_interconnect_1_uart0_s1_begintransfer;                 // mm_interconnect_1:uart0_s1_begintransfer -> uart0:begintransfer
	wire         mm_interconnect_1_uart0_s1_write;                         // mm_interconnect_1:uart0_s1_write -> uart0:write_n
	wire  [15:0] mm_interconnect_1_uart0_s1_writedata;                     // mm_interconnect_1:uart0_s1_writedata -> uart0:writedata
	wire         mm_interconnect_1_uart1_s1_chipselect;                    // mm_interconnect_1:uart1_s1_chipselect -> uart1:chipselect
	wire  [15:0] mm_interconnect_1_uart1_s1_readdata;                      // uart1:readdata -> mm_interconnect_1:uart1_s1_readdata
	wire   [2:0] mm_interconnect_1_uart1_s1_address;                       // mm_interconnect_1:uart1_s1_address -> uart1:address
	wire         mm_interconnect_1_uart1_s1_read;                          // mm_interconnect_1:uart1_s1_read -> uart1:read_n
	wire         mm_interconnect_1_uart1_s1_begintransfer;                 // mm_interconnect_1:uart1_s1_begintransfer -> uart1:begintransfer
	wire         mm_interconnect_1_uart1_s1_write;                         // mm_interconnect_1:uart1_s1_write -> uart1:write_n
	wire  [15:0] mm_interconnect_1_uart1_s1_writedata;                     // mm_interconnect_1:uart1_s1_writedata -> uart1:writedata
	wire  [31:0] mm_interconnect_1_spi_s1_readdata;                        // spi:avs_readdata -> mm_interconnect_1:spi_s1_readdata
	wire   [0:0] mm_interconnect_1_spi_s1_address;                         // mm_interconnect_1:spi_s1_address -> spi:avs_address
	wire         mm_interconnect_1_spi_s1_read;                            // mm_interconnect_1:spi_s1_read -> spi:avs_read
	wire         mm_interconnect_1_spi_s1_write;                           // mm_interconnect_1:spi_s1_write -> spi:avs_write
	wire  [31:0] mm_interconnect_1_spi_s1_writedata;                       // mm_interconnect_1:spi_s1_writedata -> spi:avs_writedata
	wire  [31:0] mm_interconnect_1_i2c_s1_readdata;                        // i2c:avs_readdata -> mm_interconnect_1:i2c_s1_readdata
	wire   [0:0] mm_interconnect_1_i2c_s1_address;                         // mm_interconnect_1:i2c_s1_address -> i2c:avs_address
	wire         mm_interconnect_1_i2c_s1_read;                            // mm_interconnect_1:i2c_s1_read -> i2c:avs_read
	wire         mm_interconnect_1_i2c_s1_write;                           // mm_interconnect_1:i2c_s1_write -> i2c:avs_write
	wire  [31:0] mm_interconnect_1_i2c_s1_writedata;                       // mm_interconnect_1:i2c_s1_writedata -> i2c:avs_writedata
	wire  [15:0] mm_interconnect_1_hostbridge_s1_readdata;                 // hostbridge:avs_readdata -> mm_interconnect_1:hostbridge_s1_readdata
	wire   [1:0] mm_interconnect_1_hostbridge_s1_address;                  // mm_interconnect_1:hostbridge_s1_address -> hostbridge:avs_address
	wire         mm_interconnect_1_hostbridge_s1_read;                     // mm_interconnect_1:hostbridge_s1_read -> hostbridge:avs_read
	wire         mm_interconnect_1_hostbridge_s1_write;                    // mm_interconnect_1:hostbridge_s1_write -> hostbridge:avs_write
	wire  [15:0] mm_interconnect_1_hostbridge_s1_writedata;                // mm_interconnect_1:hostbridge_s1_writedata -> hostbridge:avs_writedata
	wire         mm_interconnect_1_led_s1_chipselect;                      // mm_interconnect_1:led_s1_chipselect -> led:chipselect
	wire  [31:0] mm_interconnect_1_led_s1_readdata;                        // led:readdata -> mm_interconnect_1:led_s1_readdata
	wire   [1:0] mm_interconnect_1_led_s1_address;                         // mm_interconnect_1:led_s1_address -> led:address
	wire         mm_interconnect_1_led_s1_write;                           // mm_interconnect_1:led_s1_write -> led:write_n
	wire  [31:0] mm_interconnect_1_led_s1_writedata;                       // mm_interconnect_1:led_s1_writedata -> led:writedata
	wire         irq_mapper_receiver6_irq;                                 // epcs:ins_irq -> irq_mapper:receiver6_irq
	wire  [31:0] nios2_fast_irq_irq;                                       // irq_mapper:sender_irq -> nios2_fast:irq
	wire         irq_mapper_receiver0_irq;                                 // irq_synchronizer:sender_irq -> irq_mapper:receiver0_irq
	wire   [0:0] irq_synchronizer_receiver_irq;                            // systimer:irq -> irq_synchronizer:receiver_irq
	wire         irq_mapper_receiver1_irq;                                 // irq_synchronizer_001:sender_irq -> irq_mapper:receiver1_irq
	wire   [0:0] irq_synchronizer_001_receiver_irq;                        // uart0:irq -> irq_synchronizer_001:receiver_irq
	wire         irq_mapper_receiver2_irq;                                 // irq_synchronizer_002:sender_irq -> irq_mapper:receiver2_irq
	wire   [0:0] irq_synchronizer_002_receiver_irq;                        // uart1:irq -> irq_synchronizer_002:receiver_irq
	wire         irq_mapper_receiver3_irq;                                 // irq_synchronizer_003:sender_irq -> irq_mapper:receiver3_irq
	wire   [0:0] irq_synchronizer_003_receiver_irq;                        // spi:ins_irq -> irq_synchronizer_003:receiver_irq
	wire         irq_mapper_receiver4_irq;                                 // irq_synchronizer_004:sender_irq -> irq_mapper:receiver4_irq
	wire   [0:0] irq_synchronizer_004_receiver_irq;                        // i2c:ins_irq -> irq_synchronizer_004:receiver_irq
	wire         irq_mapper_receiver5_irq;                                 // irq_synchronizer_005:sender_irq -> irq_mapper:receiver5_irq
	wire   [0:0] irq_synchronizer_005_receiver_irq;                        // hostbridge:ins_irq -> irq_synchronizer_005:receiver_irq
	wire         rst_controller_reset_out_reset;                           // rst_controller:reset_out -> [rst_controller_001:reset_in0, rst_controller_002:reset_in0]
	wire         rst_controller_001_reset_out_reset;                       // rst_controller_001:reset_out -> [epcs:rsi_reset, irq_mapper:reset, irq_synchronizer:sender_reset, irq_synchronizer_001:sender_reset, irq_synchronizer_002:sender_reset, irq_synchronizer_003:sender_reset, irq_synchronizer_004:sender_reset, irq_synchronizer_005:sender_reset, mm_interconnect_0:nios2_fast_reset_reset_bridge_in_reset_reset, nios2_fast:reset_n, peripheral_bridge:s0_reset, rst_translator:in_reset, sdram:reset_n, ufm:reset_n]
	wire         rst_controller_001_reset_out_reset_req;                   // rst_controller_001:reset_req -> [nios2_fast:reset_req, rst_translator:reset_req_in]
	wire         rst_controller_002_reset_out_reset;                       // rst_controller_002:reset_out -> [chipid:reset, dual_boot_0:nreset, hostbridge:reset, i2c:rsi_reset, irq_synchronizer:receiver_reset, irq_synchronizer_001:receiver_reset, irq_synchronizer_002:receiver_reset, irq_synchronizer_003:receiver_reset, irq_synchronizer_004:receiver_reset, irq_synchronizer_005:receiver_reset, led:reset_n, mm_interconnect_1:peripheral_bridge_m0_reset_reset_bridge_in_reset_reset, peripheral_bridge:m0_reset, pfc:rsi_reset, servo:rsi_reset, spi:rsi_reset, sysid:reset_n, systimer:reset_n, uart0:reset_n, uart1:reset_n]

	altchip_id_avm_wrapper #(
		.DEVICE_FAMILY      ("MAX 10"),
		.VALIDITY_ASSERTION ("WAIT")
	) chipid (
		.clk                (clk_25m_clk),                                 //  clock.clk
		.reset              (rst_controller_002_reset_out_reset),          //  reset.reset
		.chipid_address     (mm_interconnect_1_chipid_chipid_address),     // chipid.address
		.chipid_read        (mm_interconnect_1_chipid_chipid_read),        //       .read
		.chipid_readdata    (mm_interconnect_1_chipid_chipid_readdata),    //       .readdata
		.chipid_waitrequest (mm_interconnect_1_chipid_chipid_waitrequest), //       .waitrequest
		.valid_read         (1'b0),                                        // (terminated)
		.valid_readdata     ()                                             // (terminated)
	);

	altera_dual_boot #(
		.INTENDED_DEVICE_FAMILY ("MAX 10"),
		.CONFIG_CYCLE           (9),
		.RESET_TIMER_CYCLE      (13)
	) dual_boot_0 (
		.clk                (clk_25m_clk),                                    //    clk.clk
		.nreset             (~rst_controller_002_reset_out_reset),            // nreset.reset_n
		.avmm_rcv_address   (mm_interconnect_1_dual_boot_0_avalon_address),   // avalon.address
		.avmm_rcv_read      (mm_interconnect_1_dual_boot_0_avalon_read),      //       .read
		.avmm_rcv_writedata (mm_interconnect_1_dual_boot_0_avalon_writedata), //       .writedata
		.avmm_rcv_write     (mm_interconnect_1_dual_boot_0_avalon_write),     //       .write
		.avmm_rcv_readdata  (mm_interconnect_1_dual_boot_0_avalon_readdata)   //       .readdata
	);

	peridot_csr_spi #(
		.DEFAULT_REG_BITRVS (0),
		.DEFAULT_REG_MODE   (0),
		.DEFAULT_REG_CLKDIV (255)
	) epcs (
		.csi_clk       (clk_100m_clk),                        //  clock.clk
		.rsi_reset     (rst_controller_001_reset_out_reset),  //  reset.reset
		.avs_address   (mm_interconnect_0_epcs_s1_address),   //     s1.address
		.avs_read      (mm_interconnect_0_epcs_s1_read),      //       .read
		.avs_readdata  (mm_interconnect_0_epcs_s1_readdata),  //       .readdata
		.avs_write     (mm_interconnect_0_epcs_s1_write),     //       .write
		.avs_writedata (mm_interconnect_0_epcs_s1_writedata), //       .writedata
		.ins_irq       (irq_mapper_receiver6_irq),            //    irq.irq
		.spi_ss_n      (epcs_ss_n),                           // export.ss_n
		.spi_sclk      (epcs_sclk),                           //       .sclk
		.spi_mosi      (epcs_mosi),                           //       .mosi
		.spi_miso      (epcs_miso)                            //       .miso
	);

	buffered_uart #(
		.DEVICE_FAMILY ("MAX 10"),
		.DIVIDER_BITS  (6),
		.DIVIDER_INIT  (53),
		.DIVIDER_FIXED (1),
		.RTSCTS_ENABLE (0),
		.DATA_BITS     (8),
		.RX_DEPTH_BITS (10),
		.TX_DEPTH_BITS (10)
	) hostbridge (
		.clk           (clk_25m_clk),                               // clock.clk
		.reset         (rst_controller_002_reset_out_reset),        // reset.reset
		.avs_address   (mm_interconnect_1_hostbridge_s1_address),   //    s1.address
		.avs_read      (mm_interconnect_1_hostbridge_s1_read),      //      .read
		.avs_readdata  (mm_interconnect_1_hostbridge_s1_readdata),  //      .readdata
		.avs_write     (mm_interconnect_1_hostbridge_s1_write),     //      .write
		.avs_writedata (mm_interconnect_1_hostbridge_s1_writedata), //      .writedata
		.ins_irq       (irq_synchronizer_005_receiver_irq),         //   irq.irq
		.coe_rxd       (hostuart_rxd),                              //  uart.rxd
		.coe_txd       (hostuart_txd),                              //      .txd
		.coe_rts       (),                                          // (terminated)
		.coe_cts       (1'b0)                                       // (terminated)
	);

	peridot_i2c i2c (
		.csi_clk       (clk_25m_clk),                        //  clock.clk
		.rsi_reset     (rst_controller_002_reset_out_reset), //  reset.reset
		.avs_address   (mm_interconnect_1_i2c_s1_address),   //     s1.address
		.avs_read      (mm_interconnect_1_i2c_s1_read),      //       .read
		.avs_readdata  (mm_interconnect_1_i2c_s1_readdata),  //       .readdata
		.avs_write     (mm_interconnect_1_i2c_s1_write),     //       .write
		.avs_writedata (mm_interconnect_1_i2c_s1_writedata), //       .writedata
		.ins_irq       (irq_synchronizer_004_receiver_irq),  //    irq.irq
		.i2c_scl       (i2c_scl),                            // export.scl
		.i2c_scl_oe    (i2c_scl_oe),                         //       .scl_oe
		.i2c_sda       (i2c_sda),                            //       .sda
		.i2c_sda_oe    (i2c_sda_oe)                          //       .sda_oe
	);

	olive_std_core_led led (
		.clk        (clk_25m_clk),                         //                 clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset), //               reset.reset_n
		.address    (mm_interconnect_1_led_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_led_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_led_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_led_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_led_s1_readdata),   //                    .readdata
		.out_port   (led_export)                           // external_connection.export
	);

	olive_std_core_nios2_fast nios2_fast (
		.clk                                 (clk_100m_clk),                                             //                       clk.clk
		.reset_n                             (~rst_controller_001_reset_out_reset),                      //                     reset.reset_n
		.reset_req                           (rst_controller_001_reset_out_reset_req),                   //                          .reset_req
		.d_address                           (nios2_fast_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_fast_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_fast_data_master_read),                              //                          .read
		.d_readdata                          (nios2_fast_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_fast_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_fast_data_master_write),                             //                          .write
		.d_writedata                         (nios2_fast_data_master_writedata),                         //                          .writedata
		.d_readdatavalid                     (nios2_fast_data_master_readdatavalid),                     //                          .readdatavalid
		.debug_mem_slave_debugaccess_to_roms (nios2_fast_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_fast_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_fast_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_fast_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_fast_instruction_master_waitrequest),                //                          .waitrequest
		.i_readdatavalid                     (nios2_fast_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (nios2_fast_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (),                                                         //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_fast_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_fast_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_fast_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_fast_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_fast_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_fast_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_fast_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_fast_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       (),                                                         // custom_instruction_master.readra
		.cpu_resetrequest                    (nios2_cpu_resetrequest),                                   //  cpu_resetrequest_conduit.cpu_resetrequest
		.cpu_resettaken                      (nios2_cpu_resettaken)                                      //                          .cpu_resettaken
	);

	altera_avalon_mm_clock_crossing_bridge #(
		.DATA_WIDTH          (32),
		.SYMBOL_WIDTH        (8),
		.HDL_ADDR_WIDTH      (9),
		.BURSTCOUNT_WIDTH    (1),
		.COMMAND_FIFO_DEPTH  (4),
		.RESPONSE_FIFO_DEPTH (4),
		.MASTER_SYNC_DEPTH   (2),
		.SLAVE_SYNC_DEPTH    (2)
	) peripheral_bridge (
		.m0_clk           (clk_25m_clk),                                          //   m0_clk.clk
		.m0_reset         (rst_controller_002_reset_out_reset),                   // m0_reset.reset
		.s0_clk           (clk_100m_clk),                                         //   s0_clk.clk
		.s0_reset         (rst_controller_001_reset_out_reset),                   // s0_reset.reset
		.s0_waitrequest   (mm_interconnect_0_peripheral_bridge_s0_waitrequest),   //       s0.waitrequest
		.s0_readdata      (mm_interconnect_0_peripheral_bridge_s0_readdata),      //         .readdata
		.s0_readdatavalid (mm_interconnect_0_peripheral_bridge_s0_readdatavalid), //         .readdatavalid
		.s0_burstcount    (mm_interconnect_0_peripheral_bridge_s0_burstcount),    //         .burstcount
		.s0_writedata     (mm_interconnect_0_peripheral_bridge_s0_writedata),     //         .writedata
		.s0_address       (mm_interconnect_0_peripheral_bridge_s0_address),       //         .address
		.s0_write         (mm_interconnect_0_peripheral_bridge_s0_write),         //         .write
		.s0_read          (mm_interconnect_0_peripheral_bridge_s0_read),          //         .read
		.s0_byteenable    (mm_interconnect_0_peripheral_bridge_s0_byteenable),    //         .byteenable
		.s0_debugaccess   (mm_interconnect_0_peripheral_bridge_s0_debugaccess),   //         .debugaccess
		.m0_waitrequest   (peripheral_bridge_m0_waitrequest),                     //       m0.waitrequest
		.m0_readdata      (peripheral_bridge_m0_readdata),                        //         .readdata
		.m0_readdatavalid (peripheral_bridge_m0_readdatavalid),                   //         .readdatavalid
		.m0_burstcount    (peripheral_bridge_m0_burstcount),                      //         .burstcount
		.m0_writedata     (peripheral_bridge_m0_writedata),                       //         .writedata
		.m0_address       (peripheral_bridge_m0_address),                         //         .address
		.m0_write         (peripheral_bridge_m0_write),                           //         .write
		.m0_read          (peripheral_bridge_m0_read),                            //         .read
		.m0_byteenable    (peripheral_bridge_m0_byteenable),                      //         .byteenable
		.m0_debugaccess   (peripheral_bridge_m0_debugaccess)                      //         .debugaccess
	);

	peridot_pfc_interface pfc (
		.csi_clk       (clk_25m_clk),                                  //        clock.clk
		.rsi_reset     (rst_controller_002_reset_out_reset),           //        reset.reset
		.avs_address   (mm_interconnect_1_pfc_avalon_slave_address),   // avalon_slave.address
		.avs_read      (mm_interconnect_1_pfc_avalon_slave_read),      //             .read
		.avs_readdata  (mm_interconnect_1_pfc_avalon_slave_readdata),  //             .readdata
		.avs_write     (mm_interconnect_1_pfc_avalon_slave_write),     //             .write
		.avs_writedata (mm_interconnect_1_pfc_avalon_slave_writedata), //             .writedata
		.coe_pfc_clk   (pfcif_pfc_clk),                                //       export.pfc_clk
		.coe_pfc_reset (pfcif_pfc_reset),                              //             .pfc_reset
		.coe_pfc_cmd   (pfcif_cmd),                                    //             .cmd
		.coe_pfc_resp  (pfcif_resp)                                    //             .resp
	);

	olive_std_core_sdram sdram (
		.clk            (clk_100m_clk),                             //   clk.clk
		.reset_n        (~rst_controller_001_reset_out_reset),      // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdr_addr),                                 //  wire.export
		.zs_ba          (sdr_ba),                                   //      .export
		.zs_cas_n       (sdr_cas_n),                                //      .export
		.zs_cke         (sdr_cke),                                  //      .export
		.zs_cs_n        (sdr_cs_n),                                 //      .export
		.zs_dq          (sdr_dq),                                   //      .export
		.zs_dqm         (sdr_dqm),                                  //      .export
		.zs_ras_n       (sdr_ras_n),                                //      .export
		.zs_we_n        (sdr_we_n)                                  //      .export
	);

	peridot_servo #(
		.PWM_CHANNEL (8),
		.CLOCKFREQ   (25000000)
	) servo (
		.csi_clk       (clk_25m_clk),                                    //        clock.clk
		.rsi_reset     (rst_controller_002_reset_out_reset),             //        reset.reset
		.avs_address   (mm_interconnect_1_servo_avalon_slave_address),   // avalon_slave.address
		.avs_read      (mm_interconnect_1_servo_avalon_slave_read),      //             .read
		.avs_readdata  (mm_interconnect_1_servo_avalon_slave_readdata),  //             .readdata
		.avs_write     (mm_interconnect_1_servo_avalon_slave_write),     //             .write
		.avs_writedata (mm_interconnect_1_servo_avalon_slave_writedata), //             .writedata
		.pwm_out       (servo_pwm),                                      //       export.pwm
		.dsm_out       (servo_dsm)                                       //             .dsm
	);

	peridot_csr_spi #(
		.DEFAULT_REG_BITRVS (0),
		.DEFAULT_REG_MODE   (0),
		.DEFAULT_REG_CLKDIV (255)
	) spi (
		.csi_clk       (clk_25m_clk),                        //  clock.clk
		.rsi_reset     (rst_controller_002_reset_out_reset), //  reset.reset
		.avs_address   (mm_interconnect_1_spi_s1_address),   //     s1.address
		.avs_read      (mm_interconnect_1_spi_s1_read),      //       .read
		.avs_readdata  (mm_interconnect_1_spi_s1_readdata),  //       .readdata
		.avs_write     (mm_interconnect_1_spi_s1_write),     //       .write
		.avs_writedata (mm_interconnect_1_spi_s1_writedata), //       .writedata
		.ins_irq       (irq_synchronizer_003_receiver_irq),  //    irq.irq
		.spi_ss_n      (spi_ss_n),                           // export.ss_n
		.spi_sclk      (spi_sclk),                           //       .sclk
		.spi_mosi      (spi_mosi),                           //       .mosi
		.spi_miso      (spi_miso)                            //       .miso
	);

	olive_std_core_sysid sysid (
		.clock    (clk_25m_clk),                                    //           clk.clk
		.reset_n  (~rst_controller_002_reset_out_reset),            //         reset.reset_n
		.readdata (mm_interconnect_1_sysid_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_1_sysid_control_slave_address)   //              .address
	);

	olive_std_core_systimer systimer (
		.clk        (clk_25m_clk),                              //   clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset),      // reset.reset_n
		.address    (mm_interconnect_1_systimer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_1_systimer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_1_systimer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_1_systimer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_1_systimer_s1_write),     //      .write_n
		.irq        (irq_synchronizer_receiver_irq)             //   irq.irq
	);

	olive_std_core_uart0 uart0 (
		.clk           (clk_25m_clk),                              //                 clk.clk
		.reset_n       (~rst_controller_002_reset_out_reset),      //               reset.reset_n
		.address       (mm_interconnect_1_uart0_s1_address),       //                  s1.address
		.begintransfer (mm_interconnect_1_uart0_s1_begintransfer), //                    .begintransfer
		.chipselect    (mm_interconnect_1_uart0_s1_chipselect),    //                    .chipselect
		.read_n        (~mm_interconnect_1_uart0_s1_read),         //                    .read_n
		.write_n       (~mm_interconnect_1_uart0_s1_write),        //                    .write_n
		.writedata     (mm_interconnect_1_uart0_s1_writedata),     //                    .writedata
		.readdata      (mm_interconnect_1_uart0_s1_readdata),      //                    .readdata
		.rxd           (uart0_rxd),                                // external_connection.export
		.txd           (uart0_txd),                                //                    .export
		.cts_n         (uart0_cts_n),                              //                    .export
		.rts_n         (uart0_rts_n),                              //                    .export
		.irq           (irq_synchronizer_001_receiver_irq)         //                 irq.irq
	);

	olive_std_core_uart0 uart1 (
		.clk           (clk_25m_clk),                              //                 clk.clk
		.reset_n       (~rst_controller_002_reset_out_reset),      //               reset.reset_n
		.address       (mm_interconnect_1_uart1_s1_address),       //                  s1.address
		.begintransfer (mm_interconnect_1_uart1_s1_begintransfer), //                    .begintransfer
		.chipselect    (mm_interconnect_1_uart1_s1_chipselect),    //                    .chipselect
		.read_n        (~mm_interconnect_1_uart1_s1_read),         //                    .read_n
		.write_n       (~mm_interconnect_1_uart1_s1_write),        //                    .write_n
		.writedata     (mm_interconnect_1_uart1_s1_writedata),     //                    .writedata
		.readdata      (mm_interconnect_1_uart1_s1_readdata),      //                    .readdata
		.rxd           (uart1_rxd),                                // external_connection.export
		.txd           (uart1_txd),                                //                    .export
		.cts_n         (uart1_cts_n),                              //                    .export
		.rts_n         (uart1_rts_n),                              //                    .export
		.irq           (irq_synchronizer_002_receiver_irq)         //                 irq.irq
	);

	altera_onchip_flash #(
		.INIT_FILENAME                       ("altera_onchip_flash.mif"),
		.INIT_FILENAME_SIM                   ("altera_onchip_flash.dat"),
		.DEVICE_FAMILY                       ("MAX 10"),
		.PART_NAME                           ("10M08SAE144C8G"),
		.DEVICE_ID                           ("08"),
		.SECTOR1_START_ADDR                  (0),
		.SECTOR1_END_ADDR                    (4095),
		.SECTOR2_START_ADDR                  (4096),
		.SECTOR2_END_ADDR                    (8191),
		.SECTOR3_START_ADDR                  (0),
		.SECTOR3_END_ADDR                    (0),
		.SECTOR4_START_ADDR                  (0),
		.SECTOR4_END_ADDR                    (0),
		.SECTOR5_START_ADDR                  (0),
		.SECTOR5_END_ADDR                    (0),
		.MIN_VALID_ADDR                      (0),
		.MAX_VALID_ADDR                      (8191),
		.MIN_UFM_VALID_ADDR                  (0),
		.MAX_UFM_VALID_ADDR                  (8191),
		.SECTOR1_MAP                         (1),
		.SECTOR2_MAP                         (2),
		.SECTOR3_MAP                         (0),
		.SECTOR4_MAP                         (0),
		.SECTOR5_MAP                         (0),
		.ADDR_RANGE1_END_ADDR                (8191),
		.ADDR_RANGE1_OFFSET                  (512),
		.ADDR_RANGE2_OFFSET                  (0),
		.AVMM_DATA_ADDR_WIDTH                (13),
		.AVMM_DATA_DATA_WIDTH                (32),
		.AVMM_DATA_BURSTCOUNT_WIDTH          (2),
		.SECTOR_READ_PROTECTION_MODE         (31),
		.FLASH_SEQ_READ_DATA_COUNT           (2),
		.FLASH_ADDR_ALIGNMENT_BITS           (1),
		.FLASH_READ_CYCLE_MAX_INDEX          (4),
		.FLASH_RESET_CYCLE_MAX_INDEX         (25),
		.FLASH_BUSY_TIMEOUT_CYCLE_MAX_INDEX  (120),
		.FLASH_ERASE_TIMEOUT_CYCLE_MAX_INDEX (35000000),
		.FLASH_WRITE_TIMEOUT_CYCLE_MAX_INDEX (30500),
		.PARALLEL_MODE                       (1),
		.READ_AND_WRITE_MODE                 (0),
		.WRAPPING_BURST_MODE                 (0),
		.IS_DUAL_BOOT                        ("True"),
		.IS_ERAM_SKIP                        ("True"),
		.IS_COMPRESSED_IMAGE                 ("True")
	) ufm (
		.clock                   (clk_100m_clk),                             //    clk.clk
		.reset_n                 (~rst_controller_001_reset_out_reset),      // nreset.reset_n
		.avmm_data_addr          (mm_interconnect_0_ufm_data_address),       //   data.address
		.avmm_data_read          (mm_interconnect_0_ufm_data_read),          //       .read
		.avmm_data_readdata      (mm_interconnect_0_ufm_data_readdata),      //       .readdata
		.avmm_data_waitrequest   (mm_interconnect_0_ufm_data_waitrequest),   //       .waitrequest
		.avmm_data_readdatavalid (mm_interconnect_0_ufm_data_readdatavalid), //       .readdatavalid
		.avmm_data_burstcount    (mm_interconnect_0_ufm_data_burstcount),    //       .burstcount
		.avmm_data_writedata     (32'b00000000000000000000000000000000),     // (terminated)
		.avmm_data_write         (1'b0),                                     // (terminated)
		.avmm_csr_addr           (1'b0),                                     // (terminated)
		.avmm_csr_read           (1'b0),                                     // (terminated)
		.avmm_csr_writedata      (32'b00000000000000000000000000000000),     // (terminated)
		.avmm_csr_write          (1'b0),                                     // (terminated)
		.avmm_csr_readdata       ()                                          // (terminated)
	);

	olive_std_core_mm_interconnect_0 mm_interconnect_0 (
		.core_clk_clk_clk                             (clk_100m_clk),                                             //                           core_clk_clk.clk
		.nios2_fast_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                       // nios2_fast_reset_reset_bridge_in_reset.reset
		.nios2_fast_data_master_address               (nios2_fast_data_master_address),                           //                 nios2_fast_data_master.address
		.nios2_fast_data_master_waitrequest           (nios2_fast_data_master_waitrequest),                       //                                       .waitrequest
		.nios2_fast_data_master_byteenable            (nios2_fast_data_master_byteenable),                        //                                       .byteenable
		.nios2_fast_data_master_read                  (nios2_fast_data_master_read),                              //                                       .read
		.nios2_fast_data_master_readdata              (nios2_fast_data_master_readdata),                          //                                       .readdata
		.nios2_fast_data_master_readdatavalid         (nios2_fast_data_master_readdatavalid),                     //                                       .readdatavalid
		.nios2_fast_data_master_write                 (nios2_fast_data_master_write),                             //                                       .write
		.nios2_fast_data_master_writedata             (nios2_fast_data_master_writedata),                         //                                       .writedata
		.nios2_fast_data_master_debugaccess           (nios2_fast_data_master_debugaccess),                       //                                       .debugaccess
		.nios2_fast_instruction_master_address        (nios2_fast_instruction_master_address),                    //          nios2_fast_instruction_master.address
		.nios2_fast_instruction_master_waitrequest    (nios2_fast_instruction_master_waitrequest),                //                                       .waitrequest
		.nios2_fast_instruction_master_read           (nios2_fast_instruction_master_read),                       //                                       .read
		.nios2_fast_instruction_master_readdata       (nios2_fast_instruction_master_readdata),                   //                                       .readdata
		.nios2_fast_instruction_master_readdatavalid  (nios2_fast_instruction_master_readdatavalid),              //                                       .readdatavalid
		.epcs_s1_address                              (mm_interconnect_0_epcs_s1_address),                        //                                epcs_s1.address
		.epcs_s1_write                                (mm_interconnect_0_epcs_s1_write),                          //                                       .write
		.epcs_s1_read                                 (mm_interconnect_0_epcs_s1_read),                           //                                       .read
		.epcs_s1_readdata                             (mm_interconnect_0_epcs_s1_readdata),                       //                                       .readdata
		.epcs_s1_writedata                            (mm_interconnect_0_epcs_s1_writedata),                      //                                       .writedata
		.nios2_fast_debug_mem_slave_address           (mm_interconnect_0_nios2_fast_debug_mem_slave_address),     //             nios2_fast_debug_mem_slave.address
		.nios2_fast_debug_mem_slave_write             (mm_interconnect_0_nios2_fast_debug_mem_slave_write),       //                                       .write
		.nios2_fast_debug_mem_slave_read              (mm_interconnect_0_nios2_fast_debug_mem_slave_read),        //                                       .read
		.nios2_fast_debug_mem_slave_readdata          (mm_interconnect_0_nios2_fast_debug_mem_slave_readdata),    //                                       .readdata
		.nios2_fast_debug_mem_slave_writedata         (mm_interconnect_0_nios2_fast_debug_mem_slave_writedata),   //                                       .writedata
		.nios2_fast_debug_mem_slave_byteenable        (mm_interconnect_0_nios2_fast_debug_mem_slave_byteenable),  //                                       .byteenable
		.nios2_fast_debug_mem_slave_waitrequest       (mm_interconnect_0_nios2_fast_debug_mem_slave_waitrequest), //                                       .waitrequest
		.nios2_fast_debug_mem_slave_debugaccess       (mm_interconnect_0_nios2_fast_debug_mem_slave_debugaccess), //                                       .debugaccess
		.peripheral_bridge_s0_address                 (mm_interconnect_0_peripheral_bridge_s0_address),           //                   peripheral_bridge_s0.address
		.peripheral_bridge_s0_write                   (mm_interconnect_0_peripheral_bridge_s0_write),             //                                       .write
		.peripheral_bridge_s0_read                    (mm_interconnect_0_peripheral_bridge_s0_read),              //                                       .read
		.peripheral_bridge_s0_readdata                (mm_interconnect_0_peripheral_bridge_s0_readdata),          //                                       .readdata
		.peripheral_bridge_s0_writedata               (mm_interconnect_0_peripheral_bridge_s0_writedata),         //                                       .writedata
		.peripheral_bridge_s0_burstcount              (mm_interconnect_0_peripheral_bridge_s0_burstcount),        //                                       .burstcount
		.peripheral_bridge_s0_byteenable              (mm_interconnect_0_peripheral_bridge_s0_byteenable),        //                                       .byteenable
		.peripheral_bridge_s0_readdatavalid           (mm_interconnect_0_peripheral_bridge_s0_readdatavalid),     //                                       .readdatavalid
		.peripheral_bridge_s0_waitrequest             (mm_interconnect_0_peripheral_bridge_s0_waitrequest),       //                                       .waitrequest
		.peripheral_bridge_s0_debugaccess             (mm_interconnect_0_peripheral_bridge_s0_debugaccess),       //                                       .debugaccess
		.sdram_s1_address                             (mm_interconnect_0_sdram_s1_address),                       //                               sdram_s1.address
		.sdram_s1_write                               (mm_interconnect_0_sdram_s1_write),                         //                                       .write
		.sdram_s1_read                                (mm_interconnect_0_sdram_s1_read),                          //                                       .read
		.sdram_s1_readdata                            (mm_interconnect_0_sdram_s1_readdata),                      //                                       .readdata
		.sdram_s1_writedata                           (mm_interconnect_0_sdram_s1_writedata),                     //                                       .writedata
		.sdram_s1_byteenable                          (mm_interconnect_0_sdram_s1_byteenable),                    //                                       .byteenable
		.sdram_s1_readdatavalid                       (mm_interconnect_0_sdram_s1_readdatavalid),                 //                                       .readdatavalid
		.sdram_s1_waitrequest                         (mm_interconnect_0_sdram_s1_waitrequest),                   //                                       .waitrequest
		.sdram_s1_chipselect                          (mm_interconnect_0_sdram_s1_chipselect),                    //                                       .chipselect
		.ufm_data_address                             (mm_interconnect_0_ufm_data_address),                       //                               ufm_data.address
		.ufm_data_read                                (mm_interconnect_0_ufm_data_read),                          //                                       .read
		.ufm_data_readdata                            (mm_interconnect_0_ufm_data_readdata),                      //                                       .readdata
		.ufm_data_burstcount                          (mm_interconnect_0_ufm_data_burstcount),                    //                                       .burstcount
		.ufm_data_readdatavalid                       (mm_interconnect_0_ufm_data_readdatavalid),                 //                                       .readdatavalid
		.ufm_data_waitrequest                         (mm_interconnect_0_ufm_data_waitrequest)                    //                                       .waitrequest
	);

	olive_std_core_mm_interconnect_1 mm_interconnect_1 (
		.peri_clk_clk_clk                                       (clk_25m_clk),                                    //                                     peri_clk_clk.clk
		.peripheral_bridge_m0_reset_reset_bridge_in_reset_reset (rst_controller_002_reset_out_reset),             // peripheral_bridge_m0_reset_reset_bridge_in_reset.reset
		.peripheral_bridge_m0_address                           (peripheral_bridge_m0_address),                   //                             peripheral_bridge_m0.address
		.peripheral_bridge_m0_waitrequest                       (peripheral_bridge_m0_waitrequest),               //                                                 .waitrequest
		.peripheral_bridge_m0_burstcount                        (peripheral_bridge_m0_burstcount),                //                                                 .burstcount
		.peripheral_bridge_m0_byteenable                        (peripheral_bridge_m0_byteenable),                //                                                 .byteenable
		.peripheral_bridge_m0_read                              (peripheral_bridge_m0_read),                      //                                                 .read
		.peripheral_bridge_m0_readdata                          (peripheral_bridge_m0_readdata),                  //                                                 .readdata
		.peripheral_bridge_m0_readdatavalid                     (peripheral_bridge_m0_readdatavalid),             //                                                 .readdatavalid
		.peripheral_bridge_m0_write                             (peripheral_bridge_m0_write),                     //                                                 .write
		.peripheral_bridge_m0_writedata                         (peripheral_bridge_m0_writedata),                 //                                                 .writedata
		.peripheral_bridge_m0_debugaccess                       (peripheral_bridge_m0_debugaccess),               //                                                 .debugaccess
		.chipid_chipid_address                                  (mm_interconnect_1_chipid_chipid_address),        //                                    chipid_chipid.address
		.chipid_chipid_read                                     (mm_interconnect_1_chipid_chipid_read),           //                                                 .read
		.chipid_chipid_readdata                                 (mm_interconnect_1_chipid_chipid_readdata),       //                                                 .readdata
		.chipid_chipid_waitrequest                              (mm_interconnect_1_chipid_chipid_waitrequest),    //                                                 .waitrequest
		.dual_boot_0_avalon_address                             (mm_interconnect_1_dual_boot_0_avalon_address),   //                               dual_boot_0_avalon.address
		.dual_boot_0_avalon_write                               (mm_interconnect_1_dual_boot_0_avalon_write),     //                                                 .write
		.dual_boot_0_avalon_read                                (mm_interconnect_1_dual_boot_0_avalon_read),      //                                                 .read
		.dual_boot_0_avalon_readdata                            (mm_interconnect_1_dual_boot_0_avalon_readdata),  //                                                 .readdata
		.dual_boot_0_avalon_writedata                           (mm_interconnect_1_dual_boot_0_avalon_writedata), //                                                 .writedata
		.hostbridge_s1_address                                  (mm_interconnect_1_hostbridge_s1_address),        //                                    hostbridge_s1.address
		.hostbridge_s1_write                                    (mm_interconnect_1_hostbridge_s1_write),          //                                                 .write
		.hostbridge_s1_read                                     (mm_interconnect_1_hostbridge_s1_read),           //                                                 .read
		.hostbridge_s1_readdata                                 (mm_interconnect_1_hostbridge_s1_readdata),       //                                                 .readdata
		.hostbridge_s1_writedata                                (mm_interconnect_1_hostbridge_s1_writedata),      //                                                 .writedata
		.i2c_s1_address                                         (mm_interconnect_1_i2c_s1_address),               //                                           i2c_s1.address
		.i2c_s1_write                                           (mm_interconnect_1_i2c_s1_write),                 //                                                 .write
		.i2c_s1_read                                            (mm_interconnect_1_i2c_s1_read),                  //                                                 .read
		.i2c_s1_readdata                                        (mm_interconnect_1_i2c_s1_readdata),              //                                                 .readdata
		.i2c_s1_writedata                                       (mm_interconnect_1_i2c_s1_writedata),             //                                                 .writedata
		.led_s1_address                                         (mm_interconnect_1_led_s1_address),               //                                           led_s1.address
		.led_s1_write                                           (mm_interconnect_1_led_s1_write),                 //                                                 .write
		.led_s1_readdata                                        (mm_interconnect_1_led_s1_readdata),              //                                                 .readdata
		.led_s1_writedata                                       (mm_interconnect_1_led_s1_writedata),             //                                                 .writedata
		.led_s1_chipselect                                      (mm_interconnect_1_led_s1_chipselect),            //                                                 .chipselect
		.pfc_avalon_slave_address                               (mm_interconnect_1_pfc_avalon_slave_address),     //                                 pfc_avalon_slave.address
		.pfc_avalon_slave_write                                 (mm_interconnect_1_pfc_avalon_slave_write),       //                                                 .write
		.pfc_avalon_slave_read                                  (mm_interconnect_1_pfc_avalon_slave_read),        //                                                 .read
		.pfc_avalon_slave_readdata                              (mm_interconnect_1_pfc_avalon_slave_readdata),    //                                                 .readdata
		.pfc_avalon_slave_writedata                             (mm_interconnect_1_pfc_avalon_slave_writedata),   //                                                 .writedata
		.servo_avalon_slave_address                             (mm_interconnect_1_servo_avalon_slave_address),   //                               servo_avalon_slave.address
		.servo_avalon_slave_write                               (mm_interconnect_1_servo_avalon_slave_write),     //                                                 .write
		.servo_avalon_slave_read                                (mm_interconnect_1_servo_avalon_slave_read),      //                                                 .read
		.servo_avalon_slave_readdata                            (mm_interconnect_1_servo_avalon_slave_readdata),  //                                                 .readdata
		.servo_avalon_slave_writedata                           (mm_interconnect_1_servo_avalon_slave_writedata), //                                                 .writedata
		.spi_s1_address                                         (mm_interconnect_1_spi_s1_address),               //                                           spi_s1.address
		.spi_s1_write                                           (mm_interconnect_1_spi_s1_write),                 //                                                 .write
		.spi_s1_read                                            (mm_interconnect_1_spi_s1_read),                  //                                                 .read
		.spi_s1_readdata                                        (mm_interconnect_1_spi_s1_readdata),              //                                                 .readdata
		.spi_s1_writedata                                       (mm_interconnect_1_spi_s1_writedata),             //                                                 .writedata
		.sysid_control_slave_address                            (mm_interconnect_1_sysid_control_slave_address),  //                              sysid_control_slave.address
		.sysid_control_slave_readdata                           (mm_interconnect_1_sysid_control_slave_readdata), //                                                 .readdata
		.systimer_s1_address                                    (mm_interconnect_1_systimer_s1_address),          //                                      systimer_s1.address
		.systimer_s1_write                                      (mm_interconnect_1_systimer_s1_write),            //                                                 .write
		.systimer_s1_readdata                                   (mm_interconnect_1_systimer_s1_readdata),         //                                                 .readdata
		.systimer_s1_writedata                                  (mm_interconnect_1_systimer_s1_writedata),        //                                                 .writedata
		.systimer_s1_chipselect                                 (mm_interconnect_1_systimer_s1_chipselect),       //                                                 .chipselect
		.uart0_s1_address                                       (mm_interconnect_1_uart0_s1_address),             //                                         uart0_s1.address
		.uart0_s1_write                                         (mm_interconnect_1_uart0_s1_write),               //                                                 .write
		.uart0_s1_read                                          (mm_interconnect_1_uart0_s1_read),                //                                                 .read
		.uart0_s1_readdata                                      (mm_interconnect_1_uart0_s1_readdata),            //                                                 .readdata
		.uart0_s1_writedata                                     (mm_interconnect_1_uart0_s1_writedata),           //                                                 .writedata
		.uart0_s1_begintransfer                                 (mm_interconnect_1_uart0_s1_begintransfer),       //                                                 .begintransfer
		.uart0_s1_chipselect                                    (mm_interconnect_1_uart0_s1_chipselect),          //                                                 .chipselect
		.uart1_s1_address                                       (mm_interconnect_1_uart1_s1_address),             //                                         uart1_s1.address
		.uart1_s1_write                                         (mm_interconnect_1_uart1_s1_write),               //                                                 .write
		.uart1_s1_read                                          (mm_interconnect_1_uart1_s1_read),                //                                                 .read
		.uart1_s1_readdata                                      (mm_interconnect_1_uart1_s1_readdata),            //                                                 .readdata
		.uart1_s1_writedata                                     (mm_interconnect_1_uart1_s1_writedata),           //                                                 .writedata
		.uart1_s1_begintransfer                                 (mm_interconnect_1_uart1_s1_begintransfer),       //                                                 .begintransfer
		.uart1_s1_chipselect                                    (mm_interconnect_1_uart1_s1_chipselect)           //                                                 .chipselect
	);

	olive_std_core_irq_mapper irq_mapper (
		.clk           (clk_100m_clk),                       //       clk.clk
		.reset         (rst_controller_001_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),           // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),           // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),           // receiver3.irq
		.receiver4_irq (irq_mapper_receiver4_irq),           // receiver4.irq
		.receiver5_irq (irq_mapper_receiver5_irq),           // receiver5.irq
		.receiver6_irq (irq_mapper_receiver6_irq),           // receiver6.irq
		.sender_irq    (nios2_fast_irq_irq)                  //    sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer (
		.receiver_clk   (clk_25m_clk),                        //       receiver_clk.clk
		.sender_clk     (clk_100m_clk),                       //         sender_clk.clk
		.receiver_reset (rst_controller_002_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_001_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_receiver_irq),      //           receiver.irq
		.sender_irq     (irq_mapper_receiver0_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_001 (
		.receiver_clk   (clk_25m_clk),                        //       receiver_clk.clk
		.sender_clk     (clk_100m_clk),                       //         sender_clk.clk
		.receiver_reset (rst_controller_002_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_001_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_001_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver1_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_002 (
		.receiver_clk   (clk_25m_clk),                        //       receiver_clk.clk
		.sender_clk     (clk_100m_clk),                       //         sender_clk.clk
		.receiver_reset (rst_controller_002_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_001_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_002_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver2_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_003 (
		.receiver_clk   (clk_25m_clk),                        //       receiver_clk.clk
		.sender_clk     (clk_100m_clk),                       //         sender_clk.clk
		.receiver_reset (rst_controller_002_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_001_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_003_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver3_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_004 (
		.receiver_clk   (clk_25m_clk),                        //       receiver_clk.clk
		.sender_clk     (clk_100m_clk),                       //         sender_clk.clk
		.receiver_reset (rst_controller_002_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_001_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_004_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver4_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_005 (
		.receiver_clk   (clk_25m_clk),                        //       receiver_clk.clk
		.sender_clk     (clk_100m_clk),                       //         sender_clk.clk
		.receiver_reset (rst_controller_002_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_001_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_005_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver5_irq)            //             sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (clk_100m_clk),                   //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (rst_controller_reset_out_reset),         // reset_in0.reset
		.clk            (clk_100m_clk),                           //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_001_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_in1      (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (rst_controller_reset_out_reset),     // reset_in0.reset
		.clk            (clk_25m_clk),                        //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
